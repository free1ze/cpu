
`timescale 1ns / 1ps
`include"ALUCU.sv"

module ALUCU_test();
	//too lazy to test
endmodule